VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM128_1RW1R
  CLASS BLOCK ;
  FOREIGN RAM128_1RW1R ;
  ORIGIN 0.000 0.000 ;
  SIZE 467.360 BY 552.160 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 465.360 63.960 467.360 64.560 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 465.360 106.120 467.360 106.720 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 465.360 148.280 467.360 148.880 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 465.360 190.440 467.360 191.040 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 465.360 232.600 467.360 233.200 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 465.360 274.760 467.360 275.360 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 465.360 316.920 467.360 317.520 ;
    END
  END A0[6]
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 2.000 105.360 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 2.000 173.360 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 2.000 241.360 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 2.000 309.360 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 2.000 377.360 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 2.000 445.360 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 2.000 513.360 ;
    END
  END A1[6]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 465.360 359.080 467.360 359.680 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 550.160 16.470 552.160 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 85.190 550.160 85.470 552.160 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 92.090 550.160 92.370 552.160 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 98.990 550.160 99.270 552.160 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 105.890 550.160 106.170 552.160 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 550.160 113.070 552.160 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 550.160 119.970 552.160 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 126.590 550.160 126.870 552.160 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 133.490 550.160 133.770 552.160 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 140.390 550.160 140.670 552.160 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 147.290 550.160 147.570 552.160 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 23.090 550.160 23.370 552.160 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 154.190 550.160 154.470 552.160 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 161.090 550.160 161.370 552.160 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 167.990 550.160 168.270 552.160 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 174.890 550.160 175.170 552.160 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 181.790 550.160 182.070 552.160 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 188.690 550.160 188.970 552.160 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 195.590 550.160 195.870 552.160 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 202.490 550.160 202.770 552.160 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 209.390 550.160 209.670 552.160 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 216.290 550.160 216.570 552.160 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 29.990 550.160 30.270 552.160 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 223.190 550.160 223.470 552.160 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 230.090 550.160 230.370 552.160 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 36.890 550.160 37.170 552.160 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 43.790 550.160 44.070 552.160 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 50.690 550.160 50.970 552.160 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 57.590 550.160 57.870 552.160 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 550.160 64.770 552.160 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 71.390 550.160 71.670 552.160 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 78.290 550.160 78.570 552.160 ;
    END
  END Do0[9]
  PIN Do1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 236.990 550.160 237.270 552.160 ;
    END
  END Do1[0]
  PIN Do1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 305.990 550.160 306.270 552.160 ;
    END
  END Do1[10]
  PIN Do1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 312.890 550.160 313.170 552.160 ;
    END
  END Do1[11]
  PIN Do1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 319.790 550.160 320.070 552.160 ;
    END
  END Do1[12]
  PIN Do1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 326.690 550.160 326.970 552.160 ;
    END
  END Do1[13]
  PIN Do1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 333.590 550.160 333.870 552.160 ;
    END
  END Do1[14]
  PIN Do1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 340.490 550.160 340.770 552.160 ;
    END
  END Do1[15]
  PIN Do1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 347.390 550.160 347.670 552.160 ;
    END
  END Do1[16]
  PIN Do1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 354.290 550.160 354.570 552.160 ;
    END
  END Do1[17]
  PIN Do1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 361.190 550.160 361.470 552.160 ;
    END
  END Do1[18]
  PIN Do1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 368.090 550.160 368.370 552.160 ;
    END
  END Do1[19]
  PIN Do1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 243.890 550.160 244.170 552.160 ;
    END
  END Do1[1]
  PIN Do1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 374.990 550.160 375.270 552.160 ;
    END
  END Do1[20]
  PIN Do1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 381.890 550.160 382.170 552.160 ;
    END
  END Do1[21]
  PIN Do1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 388.790 550.160 389.070 552.160 ;
    END
  END Do1[22]
  PIN Do1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 395.690 550.160 395.970 552.160 ;
    END
  END Do1[23]
  PIN Do1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 402.590 550.160 402.870 552.160 ;
    END
  END Do1[24]
  PIN Do1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 409.490 550.160 409.770 552.160 ;
    END
  END Do1[25]
  PIN Do1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 416.390 550.160 416.670 552.160 ;
    END
  END Do1[26]
  PIN Do1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 423.290 550.160 423.570 552.160 ;
    END
  END Do1[27]
  PIN Do1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 430.190 550.160 430.470 552.160 ;
    END
  END Do1[28]
  PIN Do1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 437.090 550.160 437.370 552.160 ;
    END
  END Do1[29]
  PIN Do1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 250.790 550.160 251.070 552.160 ;
    END
  END Do1[2]
  PIN Do1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 443.990 550.160 444.270 552.160 ;
    END
  END Do1[30]
  PIN Do1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 450.890 550.160 451.170 552.160 ;
    END
  END Do1[31]
  PIN Do1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 257.690 550.160 257.970 552.160 ;
    END
  END Do1[3]
  PIN Do1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 264.590 550.160 264.870 552.160 ;
    END
  END Do1[4]
  PIN Do1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 271.490 550.160 271.770 552.160 ;
    END
  END Do1[5]
  PIN Do1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 278.390 550.160 278.670 552.160 ;
    END
  END Do1[6]
  PIN Do1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 285.290 550.160 285.570 552.160 ;
    END
  END Do1[7]
  PIN Do1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 292.190 550.160 292.470 552.160 ;
    END
  END Do1[8]
  PIN Do1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 299.090 550.160 299.370 552.160 ;
    END
  END Do1[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 465.360 21.800 467.360 22.400 ;
    END
  END EN0
  PIN EN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.000 37.360 ;
    END
  END EN1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.580 2.480 23.180 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.180 2.480 176.780 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.780 2.480 330.380 549.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 549.680 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 465.360 401.240 467.360 401.840 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 465.360 443.400 467.360 444.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 465.360 485.560 467.360 486.160 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 465.360 527.720 467.360 528.320 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 2.570 2.635 464.790 549.630 ;
      LAYER li1 ;
        RECT 2.760 2.635 464.600 549.525 ;
      LAYER met1 ;
        RECT 0.070 0.040 466.830 552.120 ;
      LAYER met2 ;
        RECT 0.100 549.880 15.910 552.150 ;
        RECT 16.750 549.880 22.810 552.150 ;
        RECT 23.650 549.880 29.710 552.150 ;
        RECT 30.550 549.880 36.610 552.150 ;
        RECT 37.450 549.880 43.510 552.150 ;
        RECT 44.350 549.880 50.410 552.150 ;
        RECT 51.250 549.880 57.310 552.150 ;
        RECT 58.150 549.880 64.210 552.150 ;
        RECT 65.050 549.880 71.110 552.150 ;
        RECT 71.950 549.880 78.010 552.150 ;
        RECT 78.850 549.880 84.910 552.150 ;
        RECT 85.750 549.880 91.810 552.150 ;
        RECT 92.650 549.880 98.710 552.150 ;
        RECT 99.550 549.880 105.610 552.150 ;
        RECT 106.450 549.880 112.510 552.150 ;
        RECT 113.350 549.880 119.410 552.150 ;
        RECT 120.250 549.880 126.310 552.150 ;
        RECT 127.150 549.880 133.210 552.150 ;
        RECT 134.050 549.880 140.110 552.150 ;
        RECT 140.950 549.880 147.010 552.150 ;
        RECT 147.850 549.880 153.910 552.150 ;
        RECT 154.750 549.880 160.810 552.150 ;
        RECT 161.650 549.880 167.710 552.150 ;
        RECT 168.550 549.880 174.610 552.150 ;
        RECT 175.450 549.880 181.510 552.150 ;
        RECT 182.350 549.880 188.410 552.150 ;
        RECT 189.250 549.880 195.310 552.150 ;
        RECT 196.150 549.880 202.210 552.150 ;
        RECT 203.050 549.880 209.110 552.150 ;
        RECT 209.950 549.880 216.010 552.150 ;
        RECT 216.850 549.880 222.910 552.150 ;
        RECT 223.750 549.880 229.810 552.150 ;
        RECT 230.650 549.880 236.710 552.150 ;
        RECT 237.550 549.880 243.610 552.150 ;
        RECT 244.450 549.880 250.510 552.150 ;
        RECT 251.350 549.880 257.410 552.150 ;
        RECT 258.250 549.880 264.310 552.150 ;
        RECT 265.150 549.880 271.210 552.150 ;
        RECT 272.050 549.880 278.110 552.150 ;
        RECT 278.950 549.880 285.010 552.150 ;
        RECT 285.850 549.880 291.910 552.150 ;
        RECT 292.750 549.880 298.810 552.150 ;
        RECT 299.650 549.880 305.710 552.150 ;
        RECT 306.550 549.880 312.610 552.150 ;
        RECT 313.450 549.880 319.510 552.150 ;
        RECT 320.350 549.880 326.410 552.150 ;
        RECT 327.250 549.880 333.310 552.150 ;
        RECT 334.150 549.880 340.210 552.150 ;
        RECT 341.050 549.880 347.110 552.150 ;
        RECT 347.950 549.880 354.010 552.150 ;
        RECT 354.850 549.880 360.910 552.150 ;
        RECT 361.750 549.880 367.810 552.150 ;
        RECT 368.650 549.880 374.710 552.150 ;
        RECT 375.550 549.880 381.610 552.150 ;
        RECT 382.450 549.880 388.510 552.150 ;
        RECT 389.350 549.880 395.410 552.150 ;
        RECT 396.250 549.880 402.310 552.150 ;
        RECT 403.150 549.880 409.210 552.150 ;
        RECT 410.050 549.880 416.110 552.150 ;
        RECT 416.950 549.880 423.010 552.150 ;
        RECT 423.850 549.880 429.910 552.150 ;
        RECT 430.750 549.880 436.810 552.150 ;
        RECT 437.650 549.880 443.710 552.150 ;
        RECT 444.550 549.880 450.610 552.150 ;
        RECT 451.450 549.880 466.810 552.150 ;
        RECT 0.100 2.280 466.810 549.880 ;
        RECT 0.100 0.010 12.230 2.280 ;
        RECT 13.070 0.010 26.490 2.280 ;
        RECT 27.330 0.010 40.750 2.280 ;
        RECT 41.590 0.010 55.010 2.280 ;
        RECT 55.850 0.010 69.270 2.280 ;
        RECT 70.110 0.010 83.530 2.280 ;
        RECT 84.370 0.010 97.790 2.280 ;
        RECT 98.630 0.010 112.050 2.280 ;
        RECT 112.890 0.010 126.310 2.280 ;
        RECT 127.150 0.010 140.570 2.280 ;
        RECT 141.410 0.010 154.830 2.280 ;
        RECT 155.670 0.010 169.090 2.280 ;
        RECT 169.930 0.010 183.350 2.280 ;
        RECT 184.190 0.010 197.610 2.280 ;
        RECT 198.450 0.010 211.870 2.280 ;
        RECT 212.710 0.010 226.130 2.280 ;
        RECT 226.970 0.010 240.390 2.280 ;
        RECT 241.230 0.010 254.650 2.280 ;
        RECT 255.490 0.010 268.910 2.280 ;
        RECT 269.750 0.010 283.170 2.280 ;
        RECT 284.010 0.010 297.430 2.280 ;
        RECT 298.270 0.010 311.690 2.280 ;
        RECT 312.530 0.010 325.950 2.280 ;
        RECT 326.790 0.010 340.210 2.280 ;
        RECT 341.050 0.010 354.470 2.280 ;
        RECT 355.310 0.010 368.730 2.280 ;
        RECT 369.570 0.010 382.990 2.280 ;
        RECT 383.830 0.010 397.250 2.280 ;
        RECT 398.090 0.010 411.510 2.280 ;
        RECT 412.350 0.010 425.770 2.280 ;
        RECT 426.610 0.010 440.030 2.280 ;
        RECT 440.870 0.010 454.290 2.280 ;
        RECT 455.130 0.010 466.810 2.280 ;
      LAYER met3 ;
        RECT 0.525 528.720 466.835 551.985 ;
        RECT 0.525 527.320 464.960 528.720 ;
        RECT 0.525 513.760 466.835 527.320 ;
        RECT 2.400 512.360 466.835 513.760 ;
        RECT 0.525 486.560 466.835 512.360 ;
        RECT 0.525 485.160 464.960 486.560 ;
        RECT 0.525 445.760 466.835 485.160 ;
        RECT 2.400 444.400 466.835 445.760 ;
        RECT 2.400 444.360 464.960 444.400 ;
        RECT 0.525 443.000 464.960 444.360 ;
        RECT 0.525 402.240 466.835 443.000 ;
        RECT 0.525 400.840 464.960 402.240 ;
        RECT 0.525 377.760 466.835 400.840 ;
        RECT 2.400 376.360 466.835 377.760 ;
        RECT 0.525 360.080 466.835 376.360 ;
        RECT 0.525 358.680 464.960 360.080 ;
        RECT 0.525 317.920 466.835 358.680 ;
        RECT 0.525 316.520 464.960 317.920 ;
        RECT 0.525 309.760 466.835 316.520 ;
        RECT 2.400 308.360 466.835 309.760 ;
        RECT 0.525 275.760 466.835 308.360 ;
        RECT 0.525 274.360 464.960 275.760 ;
        RECT 0.525 241.760 466.835 274.360 ;
        RECT 2.400 240.360 466.835 241.760 ;
        RECT 0.525 233.600 466.835 240.360 ;
        RECT 0.525 232.200 464.960 233.600 ;
        RECT 0.525 191.440 466.835 232.200 ;
        RECT 0.525 190.040 464.960 191.440 ;
        RECT 0.525 173.760 466.835 190.040 ;
        RECT 2.400 172.360 466.835 173.760 ;
        RECT 0.525 149.280 466.835 172.360 ;
        RECT 0.525 147.880 464.960 149.280 ;
        RECT 0.525 107.120 466.835 147.880 ;
        RECT 0.525 105.760 464.960 107.120 ;
        RECT 2.400 105.720 464.960 105.760 ;
        RECT 2.400 104.360 466.835 105.720 ;
        RECT 0.525 64.960 466.835 104.360 ;
        RECT 0.525 63.560 464.960 64.960 ;
        RECT 0.525 37.760 466.835 63.560 ;
        RECT 2.400 36.360 466.835 37.760 ;
        RECT 0.525 22.800 466.835 36.360 ;
        RECT 0.525 21.400 464.960 22.800 ;
        RECT 0.525 0.175 466.835 21.400 ;
      LAYER met4 ;
        RECT 3.055 550.080 455.105 550.625 ;
        RECT 3.055 2.895 17.880 550.080 ;
        RECT 20.280 2.895 21.180 550.080 ;
        RECT 23.580 2.895 171.480 550.080 ;
        RECT 173.880 2.895 174.780 550.080 ;
        RECT 177.180 2.895 325.080 550.080 ;
        RECT 327.480 2.895 328.380 550.080 ;
        RECT 330.780 2.895 455.105 550.080 ;
  END
END RAM128_1RW1R
END LIBRARY

