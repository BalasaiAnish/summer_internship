VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM128_1RW1R
  CLASS BLOCK ;
  FOREIGN RAM128_1RW1R ;
  ORIGIN 0.000 0.000 ;
  SIZE 414.000 BY 552.160 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 412.000 63.960 414.000 64.560 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 412.000 106.120 414.000 106.720 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 412.000 148.280 414.000 148.880 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 412.000 190.440 414.000 191.040 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 412.000 232.600 414.000 233.200 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 412.000 274.760 414.000 275.360 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 412.000 316.920 414.000 317.520 ;
    END
  END A0[6]
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 2.000 105.360 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 2.000 173.360 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 2.000 241.360 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 2.000 309.360 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 2.000 377.360 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 2.000 445.360 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 2.000 513.360 ;
    END
  END A1[6]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 412.000 359.080 414.000 359.680 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 3.770 550.160 4.050 552.160 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 68.170 550.160 68.450 552.160 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 74.610 550.160 74.890 552.160 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 81.050 550.160 81.330 552.160 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 87.490 550.160 87.770 552.160 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 93.930 550.160 94.210 552.160 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 100.370 550.160 100.650 552.160 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 106.810 550.160 107.090 552.160 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 113.250 550.160 113.530 552.160 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 550.160 119.970 552.160 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 126.130 550.160 126.410 552.160 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 10.210 550.160 10.490 552.160 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 132.570 550.160 132.850 552.160 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 139.010 550.160 139.290 552.160 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 145.450 550.160 145.730 552.160 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 151.890 550.160 152.170 552.160 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 158.330 550.160 158.610 552.160 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 164.770 550.160 165.050 552.160 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 171.210 550.160 171.490 552.160 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 177.650 550.160 177.930 552.160 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 184.090 550.160 184.370 552.160 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 190.530 550.160 190.810 552.160 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 16.650 550.160 16.930 552.160 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 196.970 550.160 197.250 552.160 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 203.410 550.160 203.690 552.160 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 23.090 550.160 23.370 552.160 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 29.530 550.160 29.810 552.160 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 35.970 550.160 36.250 552.160 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 42.410 550.160 42.690 552.160 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 48.850 550.160 49.130 552.160 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 55.290 550.160 55.570 552.160 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 61.730 550.160 62.010 552.160 ;
    END
  END Do0[9]
  PIN Do1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 209.850 550.160 210.130 552.160 ;
    END
  END Do1[0]
  PIN Do1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 274.250 550.160 274.530 552.160 ;
    END
  END Do1[10]
  PIN Do1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 280.690 550.160 280.970 552.160 ;
    END
  END Do1[11]
  PIN Do1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 287.130 550.160 287.410 552.160 ;
    END
  END Do1[12]
  PIN Do1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 293.570 550.160 293.850 552.160 ;
    END
  END Do1[13]
  PIN Do1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 300.010 550.160 300.290 552.160 ;
    END
  END Do1[14]
  PIN Do1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 306.450 550.160 306.730 552.160 ;
    END
  END Do1[15]
  PIN Do1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 312.890 550.160 313.170 552.160 ;
    END
  END Do1[16]
  PIN Do1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 319.330 550.160 319.610 552.160 ;
    END
  END Do1[17]
  PIN Do1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 325.770 550.160 326.050 552.160 ;
    END
  END Do1[18]
  PIN Do1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 332.210 550.160 332.490 552.160 ;
    END
  END Do1[19]
  PIN Do1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 216.290 550.160 216.570 552.160 ;
    END
  END Do1[1]
  PIN Do1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 338.650 550.160 338.930 552.160 ;
    END
  END Do1[20]
  PIN Do1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 345.090 550.160 345.370 552.160 ;
    END
  END Do1[21]
  PIN Do1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 351.530 550.160 351.810 552.160 ;
    END
  END Do1[22]
  PIN Do1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 357.970 550.160 358.250 552.160 ;
    END
  END Do1[23]
  PIN Do1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 364.410 550.160 364.690 552.160 ;
    END
  END Do1[24]
  PIN Do1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 370.850 550.160 371.130 552.160 ;
    END
  END Do1[25]
  PIN Do1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 377.290 550.160 377.570 552.160 ;
    END
  END Do1[26]
  PIN Do1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 383.730 550.160 384.010 552.160 ;
    END
  END Do1[27]
  PIN Do1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 390.170 550.160 390.450 552.160 ;
    END
  END Do1[28]
  PIN Do1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 396.610 550.160 396.890 552.160 ;
    END
  END Do1[29]
  PIN Do1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 222.730 550.160 223.010 552.160 ;
    END
  END Do1[2]
  PIN Do1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 403.050 550.160 403.330 552.160 ;
    END
  END Do1[30]
  PIN Do1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 409.490 550.160 409.770 552.160 ;
    END
  END Do1[31]
  PIN Do1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 229.170 550.160 229.450 552.160 ;
    END
  END Do1[3]
  PIN Do1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 235.610 550.160 235.890 552.160 ;
    END
  END Do1[4]
  PIN Do1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 242.050 550.160 242.330 552.160 ;
    END
  END Do1[5]
  PIN Do1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 248.490 550.160 248.770 552.160 ;
    END
  END Do1[6]
  PIN Do1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 254.930 550.160 255.210 552.160 ;
    END
  END Do1[7]
  PIN Do1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 261.370 550.160 261.650 552.160 ;
    END
  END Do1[8]
  PIN Do1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 267.810 550.160 268.090 552.160 ;
    END
  END Do1[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 412.000 21.800 414.000 22.400 ;
    END
  END EN0
  PIN EN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.000 37.360 ;
    END
  END EN1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.580 2.480 23.180 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.180 2.480 176.780 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.780 2.480 330.380 549.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 549.680 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 412.000 401.240 414.000 401.840 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 412.000 443.400 414.000 444.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 412.000 485.560 414.000 486.160 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 412.000 527.720 414.000 528.320 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 2.570 2.635 411.430 549.630 ;
      LAYER li1 ;
        RECT 2.760 2.635 411.240 549.525 ;
      LAYER met1 ;
        RECT 0.070 0.040 413.470 552.120 ;
      LAYER met2 ;
        RECT 0.100 549.880 3.490 552.150 ;
        RECT 4.330 549.880 9.930 552.150 ;
        RECT 10.770 549.880 16.370 552.150 ;
        RECT 17.210 549.880 22.810 552.150 ;
        RECT 23.650 549.880 29.250 552.150 ;
        RECT 30.090 549.880 35.690 552.150 ;
        RECT 36.530 549.880 42.130 552.150 ;
        RECT 42.970 549.880 48.570 552.150 ;
        RECT 49.410 549.880 55.010 552.150 ;
        RECT 55.850 549.880 61.450 552.150 ;
        RECT 62.290 549.880 67.890 552.150 ;
        RECT 68.730 549.880 74.330 552.150 ;
        RECT 75.170 549.880 80.770 552.150 ;
        RECT 81.610 549.880 87.210 552.150 ;
        RECT 88.050 549.880 93.650 552.150 ;
        RECT 94.490 549.880 100.090 552.150 ;
        RECT 100.930 549.880 106.530 552.150 ;
        RECT 107.370 549.880 112.970 552.150 ;
        RECT 113.810 549.880 119.410 552.150 ;
        RECT 120.250 549.880 125.850 552.150 ;
        RECT 126.690 549.880 132.290 552.150 ;
        RECT 133.130 549.880 138.730 552.150 ;
        RECT 139.570 549.880 145.170 552.150 ;
        RECT 146.010 549.880 151.610 552.150 ;
        RECT 152.450 549.880 158.050 552.150 ;
        RECT 158.890 549.880 164.490 552.150 ;
        RECT 165.330 549.880 170.930 552.150 ;
        RECT 171.770 549.880 177.370 552.150 ;
        RECT 178.210 549.880 183.810 552.150 ;
        RECT 184.650 549.880 190.250 552.150 ;
        RECT 191.090 549.880 196.690 552.150 ;
        RECT 197.530 549.880 203.130 552.150 ;
        RECT 203.970 549.880 209.570 552.150 ;
        RECT 210.410 549.880 216.010 552.150 ;
        RECT 216.850 549.880 222.450 552.150 ;
        RECT 223.290 549.880 228.890 552.150 ;
        RECT 229.730 549.880 235.330 552.150 ;
        RECT 236.170 549.880 241.770 552.150 ;
        RECT 242.610 549.880 248.210 552.150 ;
        RECT 249.050 549.880 254.650 552.150 ;
        RECT 255.490 549.880 261.090 552.150 ;
        RECT 261.930 549.880 267.530 552.150 ;
        RECT 268.370 549.880 273.970 552.150 ;
        RECT 274.810 549.880 280.410 552.150 ;
        RECT 281.250 549.880 286.850 552.150 ;
        RECT 287.690 549.880 293.290 552.150 ;
        RECT 294.130 549.880 299.730 552.150 ;
        RECT 300.570 549.880 306.170 552.150 ;
        RECT 307.010 549.880 312.610 552.150 ;
        RECT 313.450 549.880 319.050 552.150 ;
        RECT 319.890 549.880 325.490 552.150 ;
        RECT 326.330 549.880 331.930 552.150 ;
        RECT 332.770 549.880 338.370 552.150 ;
        RECT 339.210 549.880 344.810 552.150 ;
        RECT 345.650 549.880 351.250 552.150 ;
        RECT 352.090 549.880 357.690 552.150 ;
        RECT 358.530 549.880 364.130 552.150 ;
        RECT 364.970 549.880 370.570 552.150 ;
        RECT 371.410 549.880 377.010 552.150 ;
        RECT 377.850 549.880 383.450 552.150 ;
        RECT 384.290 549.880 389.890 552.150 ;
        RECT 390.730 549.880 396.330 552.150 ;
        RECT 397.170 549.880 402.770 552.150 ;
        RECT 403.610 549.880 409.210 552.150 ;
        RECT 410.050 549.880 413.440 552.150 ;
        RECT 0.100 2.280 413.440 549.880 ;
        RECT 0.100 0.010 6.710 2.280 ;
        RECT 7.550 0.010 19.590 2.280 ;
        RECT 20.430 0.010 32.470 2.280 ;
        RECT 33.310 0.010 45.350 2.280 ;
        RECT 46.190 0.010 58.230 2.280 ;
        RECT 59.070 0.010 71.110 2.280 ;
        RECT 71.950 0.010 83.990 2.280 ;
        RECT 84.830 0.010 96.870 2.280 ;
        RECT 97.710 0.010 109.750 2.280 ;
        RECT 110.590 0.010 122.630 2.280 ;
        RECT 123.470 0.010 135.510 2.280 ;
        RECT 136.350 0.010 148.390 2.280 ;
        RECT 149.230 0.010 161.270 2.280 ;
        RECT 162.110 0.010 174.150 2.280 ;
        RECT 174.990 0.010 187.030 2.280 ;
        RECT 187.870 0.010 199.910 2.280 ;
        RECT 200.750 0.010 212.790 2.280 ;
        RECT 213.630 0.010 225.670 2.280 ;
        RECT 226.510 0.010 238.550 2.280 ;
        RECT 239.390 0.010 251.430 2.280 ;
        RECT 252.270 0.010 264.310 2.280 ;
        RECT 265.150 0.010 277.190 2.280 ;
        RECT 278.030 0.010 290.070 2.280 ;
        RECT 290.910 0.010 302.950 2.280 ;
        RECT 303.790 0.010 315.830 2.280 ;
        RECT 316.670 0.010 328.710 2.280 ;
        RECT 329.550 0.010 341.590 2.280 ;
        RECT 342.430 0.010 354.470 2.280 ;
        RECT 355.310 0.010 367.350 2.280 ;
        RECT 368.190 0.010 380.230 2.280 ;
        RECT 381.070 0.010 393.110 2.280 ;
        RECT 393.950 0.010 405.990 2.280 ;
        RECT 406.830 0.010 413.440 2.280 ;
      LAYER met3 ;
        RECT 0.985 528.720 413.015 551.985 ;
        RECT 0.985 527.320 411.600 528.720 ;
        RECT 0.985 513.760 413.015 527.320 ;
        RECT 2.400 512.360 413.015 513.760 ;
        RECT 0.985 486.560 413.015 512.360 ;
        RECT 0.985 485.160 411.600 486.560 ;
        RECT 0.985 445.760 413.015 485.160 ;
        RECT 2.400 444.400 413.015 445.760 ;
        RECT 2.400 444.360 411.600 444.400 ;
        RECT 0.985 443.000 411.600 444.360 ;
        RECT 0.985 402.240 413.015 443.000 ;
        RECT 0.985 400.840 411.600 402.240 ;
        RECT 0.985 377.760 413.015 400.840 ;
        RECT 2.400 376.360 413.015 377.760 ;
        RECT 0.985 360.080 413.015 376.360 ;
        RECT 0.985 358.680 411.600 360.080 ;
        RECT 0.985 317.920 413.015 358.680 ;
        RECT 0.985 316.520 411.600 317.920 ;
        RECT 0.985 309.760 413.015 316.520 ;
        RECT 2.400 308.360 413.015 309.760 ;
        RECT 0.985 275.760 413.015 308.360 ;
        RECT 0.985 274.360 411.600 275.760 ;
        RECT 0.985 241.760 413.015 274.360 ;
        RECT 2.400 240.360 413.015 241.760 ;
        RECT 0.985 233.600 413.015 240.360 ;
        RECT 0.985 232.200 411.600 233.600 ;
        RECT 0.985 191.440 413.015 232.200 ;
        RECT 0.985 190.040 411.600 191.440 ;
        RECT 0.985 173.760 413.015 190.040 ;
        RECT 2.400 172.360 413.015 173.760 ;
        RECT 0.985 149.280 413.015 172.360 ;
        RECT 0.985 147.880 411.600 149.280 ;
        RECT 0.985 107.120 413.015 147.880 ;
        RECT 0.985 105.760 411.600 107.120 ;
        RECT 2.400 105.720 411.600 105.760 ;
        RECT 2.400 104.360 413.015 105.720 ;
        RECT 0.985 64.960 413.015 104.360 ;
        RECT 0.985 63.560 411.600 64.960 ;
        RECT 0.985 37.760 413.015 63.560 ;
        RECT 2.400 36.360 413.015 37.760 ;
        RECT 0.985 22.800 413.015 36.360 ;
        RECT 0.985 21.400 411.600 22.800 ;
        RECT 0.985 0.175 413.015 21.400 ;
      LAYER met4 ;
        RECT 2.135 7.655 17.880 548.585 ;
        RECT 20.280 7.655 21.180 548.585 ;
        RECT 23.580 7.655 171.480 548.585 ;
        RECT 173.880 7.655 174.780 548.585 ;
        RECT 177.180 7.655 325.080 548.585 ;
        RECT 327.480 7.655 328.380 548.585 ;
        RECT 330.780 7.655 408.185 548.585 ;
  END
END RAM128_1RW1R
END LIBRARY

